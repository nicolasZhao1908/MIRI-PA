module sb #()();
    
endmodule
